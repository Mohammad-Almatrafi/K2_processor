module JCF_Logic (
    ZF,
    CF,
    J,
    D,
    C,
    S_reg,
    JCF,
    DataMemEn,
    Data_selector
);

  input logic J;
  input logic C, CF, ZF;
  input logic S_reg;
  input logic [1:0] D;
  output logic Data_selector, DataMemEn, JCF;

  logic inter;
  logic muxOut;
  assign muxOut = J ? ZF : CF;
  assign inter = muxOut & ((~S_reg & J) | (~S_reg & C));
  assign JCF = (J & ~C) | inter;
  assign Data_selector = J & C & S_reg;
  assign DataMemEn = S_reg & D[0] & D[1] & C;
endmodule
