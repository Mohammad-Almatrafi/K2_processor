// module register_ALU #(
//     parameter bits = 8
// );



// endmodule
